module BGU (
    
);
    
endmodule