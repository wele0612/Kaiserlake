module HCU (
);
    
endmodule